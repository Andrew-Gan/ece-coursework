module lab8-5( );


endmodule

